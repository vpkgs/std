module std
